interface operation;
  logic [3:0] a;
  logic [3:0] b;
  logic [5:0] c_out;
endinterface  
